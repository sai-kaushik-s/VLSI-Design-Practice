magic
tech scmos
timestamp 1597071209
<< nwell >>
rect -16 -4 50 12
rect 67 -4 105 12
<< polysilicon >>
rect 1 10 4 15
rect 29 10 32 15
rect 85 10 88 15
rect 1 -21 4 -2
rect 29 -21 32 -2
rect 85 -10 88 -2
rect 65 -15 88 -10
rect 85 -21 88 -15
rect 1 -38 4 -33
rect 29 -38 32 -33
rect 85 -38 88 -33
<< ndiffusion >>
rect -13 -28 1 -21
rect -13 -33 -9 -28
rect -4 -33 1 -28
rect 4 -25 29 -21
rect 4 -30 14 -25
rect 19 -30 29 -25
rect 4 -33 29 -30
rect 32 -27 47 -21
rect 32 -32 37 -27
rect 42 -32 47 -27
rect 32 -33 47 -32
rect 69 -27 85 -21
rect 69 -32 74 -27
rect 79 -32 85 -27
rect 69 -33 85 -32
rect 88 -24 103 -21
rect 88 -29 95 -24
rect 100 -29 103 -24
rect 88 -33 103 -29
<< pdiffusion >>
rect -13 9 1 10
rect -13 4 -9 9
rect -4 4 1 9
rect -13 -2 1 4
rect 4 -2 29 10
rect 32 4 47 10
rect 32 -1 37 4
rect 42 -1 47 4
rect 32 -2 47 -1
rect 69 9 85 10
rect 69 4 74 9
rect 79 4 85 9
rect 69 -2 85 4
rect 88 4 103 10
rect 88 -1 95 4
rect 100 -1 103 4
rect 88 -2 103 -1
<< metal1 >>
rect -9 18 0 23
rect 5 18 15 23
rect 20 18 35 23
rect 40 18 79 23
rect -9 9 -4 18
rect 74 9 79 18
rect 37 -10 42 -1
rect 95 -10 100 -1
rect 14 -15 60 -10
rect 95 -15 109 -10
rect 14 -25 19 -15
rect -9 -28 -4 -27
rect 95 -24 100 -15
rect -9 -41 -4 -33
rect 37 -41 42 -32
rect 74 -41 79 -32
rect -9 -46 2 -41
rect 7 -46 17 -41
rect 22 -46 41 -41
rect 46 -46 79 -41
<< ntransistor >>
rect 1 -33 4 -21
rect 29 -33 32 -21
rect 85 -33 88 -21
<< ptransistor >>
rect 1 -2 4 10
rect 29 -2 32 10
rect 85 -2 88 10
<< polycontact >>
rect 60 -15 65 -10
<< ndcontact >>
rect -9 -33 -4 -28
rect 14 -30 19 -25
rect 37 -32 42 -27
rect 74 -32 79 -27
rect 95 -29 100 -24
<< pdcontact >>
rect -9 4 -4 9
rect 37 -1 42 4
rect 74 4 79 9
rect 95 -1 100 4
<< psubstratepcontact >>
rect 2 -46 7 -41
rect 17 -46 22 -41
rect 41 -46 46 -41
<< nsubstratencontact >>
rect 0 18 5 23
rect 15 18 20 23
rect 35 18 40 23
<< labels >>
rlabel metal1 -2 20 -2 20 5 VDD!
rlabel metal1 -2 -44 -2 -44 1 GND!
rlabel polysilicon 3 -9 3 -9 1 A
rlabel polysilicon 31 -9 31 -9 1 B
rlabel metal1 107 -13 107 -13 7 Y
<< end >>
