`include "wallaceTreeMultiplier.v"

module top;

    reg [31:0] A, B;
    wire [63:0] C;

    wallaceTreeMultiplier mu(A, B, C);

    initial
    begin
        $dumpfile("wallaceTreeMultiplier_tb.vcd");
        $dumpvars(0, top);
    #5
        A = 32'b1000_0000_0000_0000_0000_0010_1000_0000;
        B = 32'b0000_0000_0000_0000_0000_0000_0110_0000;
    #5
        A = 32'b1000_0110_0000_1000_0100_0010_1001_1011;
        B = 32'b0011_1100_0110_0101_0010_1100_0110_0001;
    #5
        A = 32'b1001_0110_0110_0100_1010_0010_1000_0000;
        B = 32'b0011_0011_0010_0011_0010_0010_0110_0101;
    #5
        A = 32'b1000_0100_0010_1100_0110_0010_1010_0011;
        B = 32'b1100_1000_0010_0100_0011_0100_0110_1000;
    #5
        A = 32'b1001_1000_1010_0110_0100_0010_1100_0011;
        B = 32'b0010_0111_0000_0110_0010_0100_0110_0100;
    #5
        A = 32'b1010_1000_0011_1010_0101_1010_1010_0100;
        B = 32'b1100_0010_0100_0110_0100_1010_0110_0100;
    #5
        A = 32'b1001_0010_1000_0100_0010_0010_1000_0100;
        B = 32'b0110_0010_0100_1000_0100_0010_0110_0000;
    end

    initial
        $monitor("Multiplicand = %d Multiplier = %d Product = %d", A, B, C);

endmodule