magic
tech scmos
timestamp 1596719686
<< nwell >>
rect -5 5 24 28
<< polysilicon >>
rect 7 16 9 18
rect 7 -9 9 8
rect 7 -15 9 -13
<< ndiffusion >>
rect 6 -13 7 -9
rect 9 -13 10 -9
<< pdiffusion >>
rect 0 8 2 16
rect 6 8 7 16
rect 9 8 10 16
rect 14 8 18 16
<< metal1 >>
rect -1 20 3 24
rect 7 20 11 24
rect 15 20 19 24
rect 23 20 24 24
rect 2 16 6 20
rect 10 1 14 8
rect -5 -3 3 1
rect 10 -3 24 1
rect 10 -9 14 -3
rect 2 -18 6 -13
rect -1 -22 3 -18
rect 7 -22 11 -18
rect 15 -22 19 -18
rect 23 -22 24 -18
<< ntransistor >>
rect 7 -13 9 -9
<< ptransistor >>
rect 7 8 9 16
<< polycontact >>
rect 3 -3 7 1
<< ndcontact >>
rect 2 -13 6 -9
rect 10 -13 14 -9
<< pdcontact >>
rect 2 8 6 16
rect 10 8 14 16
<< psubstratepcontact >>
rect -5 -22 -1 -18
rect 3 -22 7 -18
rect 11 -22 15 -18
rect 19 -22 23 -18
<< nsubstratencontact >>
rect -5 20 -1 24
rect 3 20 7 24
rect 11 20 15 24
rect 19 20 23 24
<< labels >>
rlabel metal1 17 22 17 22 1 vdd!
rlabel metal1 17 -20 17 -20 1 gnd!
rlabel metal1 -5 -3 -5 1 3 vin
rlabel metal1 24 -3 24 1 7 vout
<< end >>
